module caller(a,b,c,out);
input a,b,c;
output out;
t_to_o_mux m1()